library IEEE;
library STD;
use IEEE.std_logic_1164.all;

entity and3 is
  port (
    i1 : in std_logic;
    i2 : in std_logic;
    i3 : in std_logic;
    o1 : out std_logic
  );
end and3;

architecture structural of and3 is
begin
  o1 <= i1 and i2 and i3;

end structural;
