-- Created by @(#)$CDS: vhdlin version IC23.1-64b 06/21/2023 09:20 (cpgbld16) $
-- on Fri Jan 16 11:18:55 2026


library IEEE;
library STD;
use IEEE.std_logic_1164.all;

entity dff_p is
  port (
    d : in std_logic;
    clk : in std_logic;
    q : out std_logic
  );
end dff_p;
