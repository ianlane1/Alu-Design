-- Created by @(#)$CDS: vhdlin version IC23.1-64b 06/21/2023 09:20 (cpgbld16) $
-- on Fri Jan 16 11:18:55 2026


library IEEE;
use IEEE.std_logic_1164.all;

entity or3 is

  port (
    i1   : in  std_logic;
    i2   : in  std_logic;
    i3   : in  std_logic;
    o1   : out std_logic);
end or3;
