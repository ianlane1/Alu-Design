-- Created by @(#)$CDS: vhdlin version IC23.1-64b 06/21/2023 09:20 (cpgbld16) $
-- on Fri Jan 16 11:18:55 2026


architecture structural of or4 is
begin
  o1 <= i1 or i2 or i3 or i4;

end structural;
