-- Created by @(#)$CDS: vhdlin version IC23.1-64b 06/21/2023 09:20 (cpgbld16) $
-- on Fri Jan 16 11:18:55 2026


architecture structural of counter is

component inverter
  port (
    input  : in  std_logic;
    output : out std_logic);
end component;

component dff_p
	port ( 
		d   : in  std_logic;
    	clk : in  std_logic;
        q   : out std_logic
	); 
end component;

component and2 
  port (
    i1	: in  std_logic;
	  i2	: in  std_logic;
    o1  : out std_logic);
end component;

component and3
  port (
    i1	: in  std_logic;
	  i2  : in  std_logic;
	  i3 	: in  std_logic;
    o1  : out std_logic
  );
end component;

component and4
  port (
    i1 : in std_logic;
    i2 : in std_logic;
    i3 : in std_logic;
    i4 : in std_logic;
    o1 : out std_logic
  );
end component;

component xor2
  port (
    i1	: in  std_logic;
	  i2	: in  std_logic;
    o1  : out std_logic
  );
end component;



for inv_0, inv_1 : inverter use entity work.inverter(structural);
for dff_0, dff_1, dff_2, dff_3, dff_4 : dff_p use entity work.dff_p(structural);
for xor2_0, xor2_1, xor2_2, xor2_3 : xor2 use entity work.xor2(structural);
for and2_0, and2_1, and2_2, and2_3, and2_4, and2_5 : and2 use entity work.and2(structural);
for and3_0 : and3 use entity work.and3(structural);
for and4_0 : and4 use entity work.and4(structural);

signal rst_bar, Q0_bar	: std_logic;
signal temp1 	: std_logic;
signal temp2	: std_logic_vector (1 downto 0);
signal temp3 	: std_logic_vector (1 downto 0);
signal temp4  : std_logic_vector (1 downto 0);
signal Q_temp	: std_logic_vector (4 downto 0);

begin

inv_0 : inverter port map (rst, rst_bar);

-- Bit 0 --
inv_1 : inverter port map (Q(0), Q0_bar);
and2_0: and2 port map (Q0_bar, rst_bar, Q_temp(0));
dff_0: dff_p port map (Q_temp(0), clk, Q(0));

-- Bit 1 --
xor2_0: xor2 port map (Q(0), Q(1), temp1);
and2_1: and2 port map (temp1, rst_bar, Q_temp(1));
dff_1: dff_p port map (Q_temp(1), clk, Q(1));

-- Bit 2 -- 
and2_2: and2 port map (Q(0), Q(1), temp2(0)); 
xor2_1: xor2 port map (Q(2), temp2(0), temp2(1));
and2_3: and2 port map (temp2(1), rst_bar, Q_temp(2));
dff_2: dff_p port map (Q_temp(2), clk, Q(2));

-- Bit 3 -- 
and3_0: and3 port map (Q(0), Q(1), Q(2), temp3(0));
xor2_2: xor2 port map (Q(3), temp3(0), temp3(1));
and2_4: and2 port map (temp3(1), rst_bar, Q_temp(3));
dff_3: dff_p port map (Q_temp(3), clk, Q(3));

-- Bit 4 --
and4_0: and4 port map(Q(0), Q(1), Q(2), Q(3), temp4(0));
xor2_3: xor2 port map(Q(4), temp4(0), temp4(1));
and2_5: and2 port map(temp4(1), rst_bar, Q_temp(4));
dff_4: dff_p port map(Q_temp(4), clk, Q(4));

end structural;
